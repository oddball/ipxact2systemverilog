
`define example_addr_width 3
`define example_data_width 32
