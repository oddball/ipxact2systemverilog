
`define example2_addr_width 2
`define example2_data_width 8
